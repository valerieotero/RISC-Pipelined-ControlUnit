`include "control_unit.v"

module control_unit_tb;


    control_unit UUT();
    initial begin
        
    end


endmodule