`include "PPU.v"
module PPU_tb;